library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity ouverture is
  port(
    E1,E2,E3,E4,E5,E6,E7,E8,E9 : in std_logic_vector(7 downto 0);
    RST, CLK, WE: in std_logic;
    S : out std_logic_vector(7 downto 0)
    );
end entity;

architecture ouverture_arch of ouverture is
signal R0_0, R1_0, R2_0, R3_0, R4_0, R5_0, R6_0, R7_0, R8_0 : std_logic_vector(7 downto 0);
signal R0_1, R1_1, R2_1, R3_1, R4_1, R5_1, R6_1, R7_1, R8_1 : std_logic_vector(7 downto 0);
signal ER0out : std_logic_vector(7 downto 0);
begin
    ER0: entity work.erosion(erosion_arch) port map(E1 => R0_0, E2 => R1_0, E3 => R2_0, E4 => R3_0, E5 => R4_0, E6 => R5_0, E7 => R6_0, E8 => R7_0, E9 => R8_0, S => ER0out);
    BR1: entity work.BancRegistre(BR_arch) port map (DATAIN => ER0out, RST => rst, CLK => clk, WE => we, R0 => R0_1, R1 => R1_1, R2 => R2_1, R3 => R3_1, R4 => R4_1, R5 => R5_1, R6 => R6_1, R7 => R7_1, R8 => R8_1);
    DI0: entity work.dilatation(dilatation_arch) port map(E1 => R0_1, E2 => R1_1, E3 => R2_1, E4 => R3_1, E5 => R4_1, E6 => R5_1, E7 => R6_1, E8 => R7_1, E9 => R8_1, S => S);
end architecture;
