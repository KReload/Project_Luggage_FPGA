library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity mul is
  port(
    A,N : in std_logic_vector(7 downto 0);
    S : out std_logic_vector(7 downto 0)
    );
end entity;

architecture mul_arch of mul is
begin
    
end architecture;
